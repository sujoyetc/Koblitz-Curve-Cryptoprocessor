//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:25:53 07/22/2014 
// Design Name: 
// Module Name:    sbm16 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sb16(a,b,c);

input wire [15:0]a;
input wire [15:0]b;
output wire [30:0]c;
assign c[0]=(a[0] & b[0]);
assign c[1]=(a[0] & b[1])^(a[1] & b[0]);
assign c[2]=(a[0] & b[2])^(a[1] & b[1])^(a[2] & b[0]);
assign c[3]=(a[0] & b[3])^(a[1] & b[2])^(a[2] & b[1])^(a[3] & b[0]);
assign c[4]=(a[0] & b[4])^(a[1] & b[3])^(a[2] & b[2])^(a[3] & b[1])^(a[4] & b[0]);
assign c[5]=(a[0] & b[5])^(a[1] & b[4])^(a[2] & b[3])^(a[3] & b[2])^(a[4] & b[1])^(a[5] & b[0]);
assign c[6]=(a[0] & b[6])^(a[1] & b[5])^(a[2] & b[4])^(a[3] & b[3])^(a[4] & b[2])^(a[5] & b[1])^(a[6] & b[0]);
assign c[7]=(a[0] & b[7])^(a[1] & b[6])^(a[2] & b[5])^(a[3] & b[4])^(a[4] & b[3])^(a[5] & b[2])^(a[6] & b[1])^(a[7] & b[0]);
assign c[8]=(a[0] & b[8])^(a[1] & b[7])^(a[2] & b[6])^(a[3] & b[5])^(a[4] & b[4])^(a[5] & b[3])^(a[6] & b[2])^(a[7] & b[1])^(a[8] & b[0]);
assign c[9]=(a[0] & b[9])^(a[1] & b[8])^(a[2] & b[7])^(a[3] & b[6])^(a[4] & b[5])^(a[5] & b[4])^(a[6] & b[3])^(a[7] & b[2])^(a[8] & b[1])^(a[9] & b[0]);
assign c[10]=(a[0] & b[10])^(a[1] & b[9])^(a[2] & b[8])^(a[3] & b[7])^(a[4] & b[6])^(a[5] & b[5])^(a[6] & b[4])^(a[7] & b[3])^(a[8] & b[2])^(a[9] & b[1])^(a[10] & b[0]);
assign c[11]=(a[0] & b[11])^(a[1] & b[10])^(a[2] & b[9])^(a[3] & b[8])^(a[4] & b[7])^(a[5] & b[6])^(a[6] & b[5])^(a[7] & b[4])^(a[8] & b[3])^(a[9] & b[2])^(a[10] & b[1])^(a[11] & b[0]);
assign c[12]=(a[0] & b[12])^(a[1] & b[11])^(a[2] & b[10])^(a[3] & b[9])^(a[4] & b[8])^(a[5] & b[7])^(a[6] & b[6])^(a[7] & b[5])^(a[8] & b[4])^(a[9] & b[3])^(a[10] & b[2])^(a[11] & b[1])^(a[12] & b[0]);
assign c[13]=(a[0] & b[13])^(a[1] & b[12])^(a[2] & b[11])^(a[3] & b[10])^(a[4] & b[9])^(a[5] & b[8])^(a[6] & b[7])^(a[7] & b[6])^(a[8] & b[5])^(a[9] & b[4])^(a[10] & b[3])^(a[11] & b[2])^(a[12] & b[1])^(a[13] & b[0]);
assign c[14]=(a[0] & b[14])^(a[1] & b[13])^(a[2] & b[12])^(a[3] & b[11])^(a[4] & b[10])^(a[5] & b[9])^(a[6] & b[8])^(a[7] & b[7])^(a[8] & b[6])^(a[9] & b[5])^(a[10] & b[4])^(a[11] & b[3])^(a[12] & b[2])^(a[13] & b[1])^(a[14] & b[0]);
assign c[15]=(a[0] & b[15])^(a[1] & b[14])^(a[2] & b[13])^(a[3] & b[12])^(a[4] & b[11])^(a[5] & b[10])^(a[6] & b[9])^(a[7] & b[8])^(a[8] & b[7])^(a[9] & b[6])^(a[10] & b[5])^(a[11] & b[4])^(a[12] & b[3])^(a[13] & b[2])^(a[14] & b[1])^(a[15] & b[0]);
assign c[16]=(a[1] & b[15])^(a[2] & b[14])^(a[3] & b[13])^(a[4] & b[12])^(a[5] & b[11])^(a[6] & b[10])^(a[7] & b[9])^(a[8] & b[8])^(a[9] & b[7])^(a[10] & b[6])^(a[11] & b[5])^(a[12] & b[4])^(a[13] & b[3])^(a[14] & b[2])^(a[15] & b[1]);
assign c[17]=(a[2] & b[15])^(a[3] & b[14])^(a[4] & b[13])^(a[5] & b[12])^(a[6] & b[11])^(a[7] & b[10])^(a[8] & b[9])^(a[9] & b[8])^(a[10] & b[7])^(a[11] & b[6])^(a[12] & b[5])^(a[13] & b[4])^(a[14] & b[3])^(a[15] & b[2]);
assign c[18]=(a[3] & b[15])^(a[4] & b[14])^(a[5] & b[13])^(a[6] & b[12])^(a[7] & b[11])^(a[8] & b[10])^(a[9] & b[9])^(a[10] & b[8])^(a[11] & b[7])^(a[12] & b[6])^(a[13] & b[5])^(a[14] & b[4])^(a[15] & b[3]);
assign c[19]=(a[4] & b[15])^(a[5] & b[14])^(a[6] & b[13])^(a[7] & b[12])^(a[8] & b[11])^(a[9] & b[10])^(a[10] & b[9])^(a[11] & b[8])^(a[12] & b[7])^(a[13] & b[6])^(a[14] & b[5])^(a[15] & b[4]);
assign c[20]=(a[5] & b[15])^(a[6] & b[14])^(a[7] & b[13])^(a[8] & b[12])^(a[9] & b[11])^(a[10] & b[10])^(a[11] & b[9])^(a[12] & b[8])^(a[13] & b[7])^(a[14] & b[6])^(a[15] & b[5]);
assign c[21]=(a[6] & b[15])^(a[7] & b[14])^(a[8] & b[13])^(a[9] & b[12])^(a[10] & b[11])^(a[11] & b[10])^(a[12] & b[9])^(a[13] & b[8])^(a[14] & b[7])^(a[15] & b[6]);
assign c[22]=(a[7] & b[15])^(a[8] & b[14])^(a[9] & b[13])^(a[10] & b[12])^(a[11] & b[11])^(a[12] & b[10])^(a[13] & b[9])^(a[14] & b[8])^(a[15] & b[7]);
assign c[23]=(a[8] & b[15])^(a[9] & b[14])^(a[10] & b[13])^(a[11] & b[12])^(a[12] & b[11])^(a[13] & b[10])^(a[14] & b[9])^(a[15] & b[8]);
assign c[24]=(a[9] & b[15])^(a[10] & b[14])^(a[11] & b[13])^(a[12] & b[12])^(a[13] & b[11])^(a[14] & b[10])^(a[15] & b[9]);
assign c[25]=(a[10] & b[15])^(a[11] & b[14])^(a[12] & b[13])^(a[13] & b[12])^(a[14] & b[11])^(a[15] & b[10]);
assign c[26]=(a[11] & b[15])^(a[12] & b[14])^(a[13] & b[13])^(a[14] & b[12])^(a[15] & b[11]);
assign c[27]=(a[12] & b[15])^(a[13] & b[14])^(a[14] & b[13])^(a[15] & b[12]);
assign c[28]=(a[13] & b[15])^(a[14] & b[14])^(a[15] & b[13]);
assign c[29]=(a[14] & b[15])^(a[15] & b[14]);
assign c[30]=(a[15] & b[15]);
endmodule
